module InstructionMemory(
	input [7:0] address,
	output reg [7:0] data
	);
	
	reg [7:0] instruction_data [0:255];

	


endmodule