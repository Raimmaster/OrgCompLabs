module InstructionMemory(
	input [7:0] address,
	output reg [7:0] instruction
	);
	
	

endmodule