module MIPS_Processor(
	input clk
	
	);

endmodule