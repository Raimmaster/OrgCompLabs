module DataMemory(
	input [1:0] address,
	input [7:0] write_data,
	input data_we,
	output [7:0] read_data
	);

	

endmodule